--******************************************************--
--        PONTIFICIA UNIVERSIDAD JAVERIANA              --
--                Disegno Digital                       --
--          Seccion de Tecnicas Digitales               --
-- 													              --
-- Titulo :                                             --
-- Fecha  :  	D:XX M:XX Y:20XX                         --
--******************************************************--
-- 													              --
-------------- Package: MyGraphs.vhd -----------------
-- 													              --
--******************************************************--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

USE WORK.MyGamePackage.ALL;

PACKAGE MyGraphs IS

CONSTANT SF : INTEGER := ShipSizeY;
CONSTANT SC : INTEGER := ShipSizeX;
CONSTANT BF : INTEGER := BulletSizeY;
CONSTANT BC : INTEGER := BulletSizeX;
CONSTANT NF : INTEGER := ScoreSizeY;
CONSTANT NC : INTEGER := ScoreSizeX;

--**************************************************************************************************--
-- 
-- Definition 
--
--**************************************************************************************************--

TYPE Matrix IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_logic_vector(7 DOWNTO 0);

--**************************************************************************************************--
-- 
-- Definition of Ship 1 figure
--
--**************************************************************************************************--

CONSTANT FigureShip1R : Matrix(0 TO SF, 0 TO SC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A8",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"A8",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"FF",	x"A8",	x"A8",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A8",	x"A8",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A8",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A8",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A8",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"A8",	x"A8",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A8",	x"A8",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF"),
(x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"A8",	x"A8",	x"A8",	x"A8",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"A8",	x"A8",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"A8",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"A8",	x"A8",	x"A8",	x"CC",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A8",	x"A8",	x"A8",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"00",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"A8",	x"A8",	x"A8",	x"A6",	x"A6",	x"A6",	x"A8",	x"A8",	x"A6",	x"A6",	x"A6",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"FF",	x"CC",	x"CC",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"CC",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"CC",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"CC",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"A8",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureShip1G : Matrix(0 TO SF, 0 TO SC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF"),
(x"00",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00"),
(x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureShip1B : Matrix(0 TO SF, 0 TO SC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66"),
(x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"00",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"00",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF"),
(x"66",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66"),
(x"66",	x"66",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Ship 2 figure
--
--**************************************************************************************************--

CONSTANT FigureShip2R : Matrix(0 TO SF, 0 TO SC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF"),
(x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6"),
(x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6"),
(x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"66",	x"66",	x"66",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"A6",	x"A6",	x"A6",	x"66",	x"66",	x"A6",	x"A6",	x"A6",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"FF",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureShip2G : Matrix(0 TO SF, 0 TO SC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6"),
(x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6"),
(x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"00"),
(x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureShip2B : Matrix(0 TO SF, 0 TO SC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"FF",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66"),
(x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"FF",	x"99",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66"),
(x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"00",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"00",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"A6"),
(x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"A6",	x"A6"),
(x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"FF",	x"99",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"66",	x"66",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"66"),
(x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"66",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"99",	x"66",	x"66",	x"66",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"00",	x"00",	x"00",	x"99",	x"99",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"A6",	x"A6",	x"A6",	x"66",	x"66",	x"A6",	x"A6",	x"A6",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"A6",	x"FF",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"A6",	x"A6",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"99",	x"FF",	x"FF",	x"00",	x"00",	x"A6",	x"A6",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"FF",	x"00",	x"A6",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"FF",	x"FF",	x"00",	x"A6",	x"A6",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"99",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

--**************************************************************************************************--
-- 
-- Definition of Bullet figure
--
--**************************************************************************************************--

CONSTANT FigureBulletR : Matrix(0 TO BF, 0 TO BC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"FF",	x"FF"),
(x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA"),
(x"FF",	x"FF",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureBulletG : Matrix(0 TO BF, 0 TO BC) := (
(x"00",	x"00",	x"00",	x"00",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"00",	x"00"),
(x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA"),
(x"00",	x"00",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureBulletB : Matrix(0 TO BF, 0 TO BC) := (
(x"66",	x"66",	x"66",	x"66",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"66",	x"66"),
(x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA"),
(x"66",	x"66",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"AA",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 0 figure
--
--**************************************************************************************************--

CONSTANT FigureNum0R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum0G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum0B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 1 figure
--
--**************************************************************************************************--

CONSTANT FigureNum1R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum1G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum1B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 2 figure
--
--**************************************************************************************************--

CONSTANT FigureNum2R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum2G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum2B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 3 figure
--
--**************************************************************************************************--

CONSTANT FigureNum3R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum3G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum3B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 4 figure
--
--**************************************************************************************************--

CONSTANT FigureNum4R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum4G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum4B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 5 figure
--
--**************************************************************************************************--

CONSTANT FigureNum5R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum5G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum5B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 6 figure
--
--**************************************************************************************************--

CONSTANT FigureNum6R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum6G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum6B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 7 figure
--
--**************************************************************************************************--

CONSTANT FigureNum7R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum7G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum7B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 8 figure
--
--**************************************************************************************************--

CONSTANT FigureNum8R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum8G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum8B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

--**************************************************************************************************--
-- 
-- Definition of Number 9 figure
--
--**************************************************************************************************--

CONSTANT FigureNum9R : Matrix(0 TO NF, 0 TO NC) := (
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"),
(x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF",	x"FF"));

CONSTANT FigureNum9G : Matrix(0 TO NF, 0 TO NC) := (
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"D7",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"),
(x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00"));

CONSTANT FigureNum9B : Matrix(0 TO NF, 0 TO NC) := (
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"00",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"),
(x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66",	x"66"));

END PACKAGE MyGraphs;

PACKAGE BODY MyGraphs IS



END MyGraphs;